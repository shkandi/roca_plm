LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

package roca_src is

type arr_26 is array(0 to 25) of std_logic_vector(7 downto 0);
type arr_256 is array (0 to 255) of std_logic_vector (7 downto 0);

end roca_src;

package body roca_src is 

end roca_src;